library verilog;
use verilog.vl_types.all;
entity tick_counter_vlg_vec_tst is
end tick_counter_vlg_vec_tst;
