library verilog;
use verilog.vl_types.all;
entity lab3ex_vlg_vec_tst is
end lab3ex_vlg_vec_tst;
